//////////////////////////DR SERAG //////////////////
////////////////Outhers:Isalm_Akram_Osama///////////

module nand_gate  (
input wire a,b,
output c
);

assign c=!(a&b);
 
endmodule

