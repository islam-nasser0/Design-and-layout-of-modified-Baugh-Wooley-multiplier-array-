//////////////////////////DR SERAG //////////////////
////////////////Outhers:Isalm_Akram_Osama///////////

module and_gate  (
input wire a,b,
output c
);

assign c=a&b;
 
endmodule